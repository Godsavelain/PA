module Decode(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_pc,
  input  [31:0] io_in_bits_inst,
  input         io_in_bits_inst_valid,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_valid,
  output [31:0] io_out_bits_pc,
  output [31:0] io_out_bits_inst,
  output [2:0]  io_out_bits_fu_code,
  output [3:0]  io_out_bits_alu_code,
  output [3:0]  io_out_bits_jmp_code,
  output [1:0]  io_out_bits_mem_code,
  output [1:0]  io_out_bits_mem_size,
  output [2:0]  io_out_bits_csr_code,
  output        io_out_bits_w_type,
  output [2:0]  io_out_bits_rs1_src,
  output [2:0]  io_out_bits_rs2_src,
  output [4:0]  io_out_bits_rs1_addr,
  output [4:0]  io_out_bits_rs2_addr,
  output [4:0]  io_out_bits_rd_addr,
  output        io_out_bits_rd_en,
  output [31:0] io_out_bits_imm,
  input         io_id_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] inst; // @[Decode.scala 15:22]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _ctrl_T = inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _ctrl_T_1 = 32'h37 == _ctrl_T; // @[Lookup.scala 31:38]
  wire  _ctrl_T_3 = 32'h17 == _ctrl_T; // @[Lookup.scala 31:38]
  wire  _ctrl_T_5 = 32'h6f == _ctrl_T; // @[Lookup.scala 31:38]
  wire [31:0] _ctrl_T_6 = inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _ctrl_T_7 = 32'h67 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_9 = 32'h63 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_11 = 32'h1063 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_13 = 32'h4063 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_15 = 32'h5063 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_17 = 32'h6063 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_19 = 32'h7063 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_21 = 32'h3 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_23 = 32'h1003 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_25 = 32'h2003 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_27 = 32'h4003 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_29 = 32'h5003 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_31 = 32'h23 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_33 = 32'h1023 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_35 = 32'h2023 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_37 = 32'h13 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_39 = 32'h2013 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_41 = 32'h3013 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_43 = 32'h4013 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_45 = 32'h6013 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_47 = 32'h7013 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire [31:0] _ctrl_T_48 = inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _ctrl_T_49 = 32'h1013 == _ctrl_T_48; // @[Lookup.scala 31:38]
  wire  _ctrl_T_51 = 32'h5013 == _ctrl_T_48; // @[Lookup.scala 31:38]
  wire  _ctrl_T_53 = 32'h40005013 == _ctrl_T_48; // @[Lookup.scala 31:38]
  wire [31:0] _ctrl_T_54 = inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _ctrl_T_55 = 32'h33 == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_57 = 32'h40000033 == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_59 = 32'h1033 == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_61 = 32'h2033 == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_63 = 32'h3033 == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_65 = 32'h4033 == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_67 = 32'h5033 == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_69 = 32'h40005033 == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_71 = 32'h6033 == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_73 = 32'h7033 == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_75 = 32'h73 == inst; // @[Lookup.scala 31:38]
  wire  _ctrl_T_77 = 32'h30200073 == inst; // @[Lookup.scala 31:38]
  wire  _ctrl_T_79 = 32'h10500073 == inst; // @[Lookup.scala 31:38]
  wire  _ctrl_T_81 = 32'h6003 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_83 = 32'h3003 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_85 = 32'h3023 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_87 = 32'h1b == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_89 = 32'h101b == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_91 = 32'h501b == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_93 = 32'h4000501b == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_95 = 32'h3b == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_97 = 32'h4000003b == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_99 = 32'h103b == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_101 = 32'h503b == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_103 = 32'h4000503b == _ctrl_T_54; // @[Lookup.scala 31:38]
  wire  _ctrl_T_105 = 32'h1073 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_107 = 32'h2073 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_109 = 32'h3073 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_111 = 32'h5073 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_113 = 32'h6073 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire  _ctrl_T_115 = 32'h7073 == _ctrl_T_6; // @[Lookup.scala 31:38]
  wire [2:0] _ctrl_T_181 = _ctrl_T_115 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_182 = _ctrl_T_113 ? 3'h4 : _ctrl_T_181; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_183 = _ctrl_T_111 ? 3'h4 : _ctrl_T_182; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_184 = _ctrl_T_109 ? 3'h4 : _ctrl_T_183; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_185 = _ctrl_T_107 ? 3'h4 : _ctrl_T_184; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_186 = _ctrl_T_105 ? 3'h4 : _ctrl_T_185; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_187 = _ctrl_T_103 ? 3'h1 : _ctrl_T_186; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_188 = _ctrl_T_101 ? 3'h1 : _ctrl_T_187; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_189 = _ctrl_T_99 ? 3'h1 : _ctrl_T_188; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_190 = _ctrl_T_97 ? 3'h1 : _ctrl_T_189; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_191 = _ctrl_T_95 ? 3'h1 : _ctrl_T_190; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_192 = _ctrl_T_93 ? 3'h1 : _ctrl_T_191; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_193 = _ctrl_T_91 ? 3'h1 : _ctrl_T_192; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_194 = _ctrl_T_89 ? 3'h1 : _ctrl_T_193; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_195 = _ctrl_T_87 ? 3'h1 : _ctrl_T_194; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_196 = _ctrl_T_85 ? 3'h3 : _ctrl_T_195; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_197 = _ctrl_T_83 ? 3'h3 : _ctrl_T_196; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_198 = _ctrl_T_81 ? 3'h3 : _ctrl_T_197; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_199 = _ctrl_T_79 ? 3'h1 : _ctrl_T_198; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_200 = _ctrl_T_77 ? 3'h4 : _ctrl_T_199; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_201 = _ctrl_T_75 ? 3'h4 : _ctrl_T_200; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_202 = _ctrl_T_73 ? 3'h1 : _ctrl_T_201; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_203 = _ctrl_T_71 ? 3'h1 : _ctrl_T_202; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_204 = _ctrl_T_69 ? 3'h1 : _ctrl_T_203; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_205 = _ctrl_T_67 ? 3'h1 : _ctrl_T_204; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_206 = _ctrl_T_65 ? 3'h1 : _ctrl_T_205; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_207 = _ctrl_T_63 ? 3'h1 : _ctrl_T_206; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_208 = _ctrl_T_61 ? 3'h1 : _ctrl_T_207; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_209 = _ctrl_T_59 ? 3'h1 : _ctrl_T_208; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_210 = _ctrl_T_57 ? 3'h1 : _ctrl_T_209; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_211 = _ctrl_T_55 ? 3'h1 : _ctrl_T_210; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_212 = _ctrl_T_53 ? 3'h1 : _ctrl_T_211; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_213 = _ctrl_T_51 ? 3'h1 : _ctrl_T_212; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_214 = _ctrl_T_49 ? 3'h1 : _ctrl_T_213; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_215 = _ctrl_T_47 ? 3'h1 : _ctrl_T_214; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_216 = _ctrl_T_45 ? 3'h1 : _ctrl_T_215; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_217 = _ctrl_T_43 ? 3'h1 : _ctrl_T_216; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_218 = _ctrl_T_41 ? 3'h1 : _ctrl_T_217; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_219 = _ctrl_T_39 ? 3'h1 : _ctrl_T_218; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_220 = _ctrl_T_37 ? 3'h1 : _ctrl_T_219; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_221 = _ctrl_T_35 ? 3'h3 : _ctrl_T_220; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_222 = _ctrl_T_33 ? 3'h3 : _ctrl_T_221; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_223 = _ctrl_T_31 ? 3'h3 : _ctrl_T_222; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_224 = _ctrl_T_29 ? 3'h3 : _ctrl_T_223; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_225 = _ctrl_T_27 ? 3'h3 : _ctrl_T_224; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_226 = _ctrl_T_25 ? 3'h3 : _ctrl_T_225; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_227 = _ctrl_T_23 ? 3'h3 : _ctrl_T_226; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_228 = _ctrl_T_21 ? 3'h3 : _ctrl_T_227; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_229 = _ctrl_T_19 ? 3'h2 : _ctrl_T_228; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_230 = _ctrl_T_17 ? 3'h2 : _ctrl_T_229; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_231 = _ctrl_T_15 ? 3'h2 : _ctrl_T_230; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_232 = _ctrl_T_13 ? 3'h2 : _ctrl_T_231; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_233 = _ctrl_T_11 ? 3'h2 : _ctrl_T_232; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_234 = _ctrl_T_9 ? 3'h2 : _ctrl_T_233; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_235 = _ctrl_T_7 ? 3'h2 : _ctrl_T_234; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_236 = _ctrl_T_5 ? 3'h2 : _ctrl_T_235; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_237 = _ctrl_T_3 ? 3'h1 : _ctrl_T_236; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_246 = _ctrl_T_103 ? 4'ha : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_247 = _ctrl_T_101 ? 4'h9 : _ctrl_T_246; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_248 = _ctrl_T_99 ? 4'h8 : _ctrl_T_247; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_249 = _ctrl_T_97 ? 4'h2 : _ctrl_T_248; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_250 = _ctrl_T_95 ? 4'h1 : _ctrl_T_249; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_251 = _ctrl_T_93 ? 4'ha : _ctrl_T_250; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_252 = _ctrl_T_91 ? 4'h9 : _ctrl_T_251; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_253 = _ctrl_T_89 ? 4'h8 : _ctrl_T_252; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_254 = _ctrl_T_87 ? 4'h1 : _ctrl_T_253; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_255 = _ctrl_T_85 ? 4'h0 : _ctrl_T_254; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_256 = _ctrl_T_83 ? 4'h0 : _ctrl_T_255; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_257 = _ctrl_T_81 ? 4'h0 : _ctrl_T_256; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_258 = _ctrl_T_79 ? 4'h0 : _ctrl_T_257; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_259 = _ctrl_T_77 ? 4'h0 : _ctrl_T_258; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_260 = _ctrl_T_75 ? 4'h0 : _ctrl_T_259; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_261 = _ctrl_T_73 ? 4'h7 : _ctrl_T_260; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_262 = _ctrl_T_71 ? 4'h6 : _ctrl_T_261; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_263 = _ctrl_T_69 ? 4'ha : _ctrl_T_262; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_264 = _ctrl_T_67 ? 4'h9 : _ctrl_T_263; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_265 = _ctrl_T_65 ? 4'h5 : _ctrl_T_264; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_266 = _ctrl_T_63 ? 4'h4 : _ctrl_T_265; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_267 = _ctrl_T_61 ? 4'h3 : _ctrl_T_266; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_268 = _ctrl_T_59 ? 4'h8 : _ctrl_T_267; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_269 = _ctrl_T_57 ? 4'h2 : _ctrl_T_268; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_270 = _ctrl_T_55 ? 4'h1 : _ctrl_T_269; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_271 = _ctrl_T_53 ? 4'ha : _ctrl_T_270; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_272 = _ctrl_T_51 ? 4'h9 : _ctrl_T_271; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_273 = _ctrl_T_49 ? 4'h8 : _ctrl_T_272; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_274 = _ctrl_T_47 ? 4'h7 : _ctrl_T_273; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_275 = _ctrl_T_45 ? 4'h6 : _ctrl_T_274; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_276 = _ctrl_T_43 ? 4'h5 : _ctrl_T_275; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_277 = _ctrl_T_41 ? 4'h4 : _ctrl_T_276; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_278 = _ctrl_T_39 ? 4'h3 : _ctrl_T_277; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_279 = _ctrl_T_37 ? 4'h1 : _ctrl_T_278; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_280 = _ctrl_T_35 ? 4'h0 : _ctrl_T_279; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_281 = _ctrl_T_33 ? 4'h0 : _ctrl_T_280; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_282 = _ctrl_T_31 ? 4'h0 : _ctrl_T_281; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_283 = _ctrl_T_29 ? 4'h0 : _ctrl_T_282; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_284 = _ctrl_T_27 ? 4'h0 : _ctrl_T_283; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_285 = _ctrl_T_25 ? 4'h0 : _ctrl_T_284; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_286 = _ctrl_T_23 ? 4'h0 : _ctrl_T_285; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_287 = _ctrl_T_21 ? 4'h0 : _ctrl_T_286; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_288 = _ctrl_T_19 ? 4'h0 : _ctrl_T_287; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_289 = _ctrl_T_17 ? 4'h0 : _ctrl_T_288; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_290 = _ctrl_T_15 ? 4'h0 : _ctrl_T_289; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_291 = _ctrl_T_13 ? 4'h0 : _ctrl_T_290; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_292 = _ctrl_T_11 ? 4'h0 : _ctrl_T_291; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_293 = _ctrl_T_9 ? 4'h0 : _ctrl_T_292; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_294 = _ctrl_T_7 ? 4'h0 : _ctrl_T_293; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_295 = _ctrl_T_5 ? 4'h0 : _ctrl_T_294; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_296 = _ctrl_T_3 ? 4'h1 : _ctrl_T_295; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_347 = _ctrl_T_19 ? 4'h8 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_348 = _ctrl_T_17 ? 4'h7 : _ctrl_T_347; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_349 = _ctrl_T_15 ? 4'h6 : _ctrl_T_348; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_350 = _ctrl_T_13 ? 4'h5 : _ctrl_T_349; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_351 = _ctrl_T_11 ? 4'h4 : _ctrl_T_350; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_352 = _ctrl_T_9 ? 4'h3 : _ctrl_T_351; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_353 = _ctrl_T_7 ? 4'h2 : _ctrl_T_352; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_354 = _ctrl_T_5 ? 4'h1 : _ctrl_T_353; // @[Lookup.scala 33:37]
  wire [3:0] _ctrl_T_355 = _ctrl_T_3 ? 4'h0 : _ctrl_T_354; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_373 = _ctrl_T_85 ? 2'h3 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_374 = _ctrl_T_83 ? 2'h2 : _ctrl_T_373; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_375 = _ctrl_T_81 ? 2'h2 : _ctrl_T_374; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_376 = _ctrl_T_79 ? 2'h0 : _ctrl_T_375; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_377 = _ctrl_T_77 ? 2'h0 : _ctrl_T_376; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_378 = _ctrl_T_75 ? 2'h0 : _ctrl_T_377; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_379 = _ctrl_T_73 ? 2'h0 : _ctrl_T_378; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_380 = _ctrl_T_71 ? 2'h0 : _ctrl_T_379; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_381 = _ctrl_T_69 ? 2'h0 : _ctrl_T_380; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_382 = _ctrl_T_67 ? 2'h0 : _ctrl_T_381; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_383 = _ctrl_T_65 ? 2'h0 : _ctrl_T_382; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_384 = _ctrl_T_63 ? 2'h0 : _ctrl_T_383; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_385 = _ctrl_T_61 ? 2'h0 : _ctrl_T_384; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_386 = _ctrl_T_59 ? 2'h0 : _ctrl_T_385; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_387 = _ctrl_T_57 ? 2'h0 : _ctrl_T_386; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_388 = _ctrl_T_55 ? 2'h0 : _ctrl_T_387; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_389 = _ctrl_T_53 ? 2'h0 : _ctrl_T_388; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_390 = _ctrl_T_51 ? 2'h0 : _ctrl_T_389; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_391 = _ctrl_T_49 ? 2'h0 : _ctrl_T_390; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_392 = _ctrl_T_47 ? 2'h0 : _ctrl_T_391; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_393 = _ctrl_T_45 ? 2'h0 : _ctrl_T_392; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_394 = _ctrl_T_43 ? 2'h0 : _ctrl_T_393; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_395 = _ctrl_T_41 ? 2'h0 : _ctrl_T_394; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_396 = _ctrl_T_39 ? 2'h0 : _ctrl_T_395; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_397 = _ctrl_T_37 ? 2'h0 : _ctrl_T_396; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_398 = _ctrl_T_35 ? 2'h3 : _ctrl_T_397; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_399 = _ctrl_T_33 ? 2'h3 : _ctrl_T_398; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_400 = _ctrl_T_31 ? 2'h3 : _ctrl_T_399; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_401 = _ctrl_T_29 ? 2'h2 : _ctrl_T_400; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_402 = _ctrl_T_27 ? 2'h2 : _ctrl_T_401; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_403 = _ctrl_T_25 ? 2'h1 : _ctrl_T_402; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_404 = _ctrl_T_23 ? 2'h1 : _ctrl_T_403; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_405 = _ctrl_T_21 ? 2'h1 : _ctrl_T_404; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_406 = _ctrl_T_19 ? 2'h0 : _ctrl_T_405; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_407 = _ctrl_T_17 ? 2'h0 : _ctrl_T_406; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_408 = _ctrl_T_15 ? 2'h0 : _ctrl_T_407; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_409 = _ctrl_T_13 ? 2'h0 : _ctrl_T_408; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_410 = _ctrl_T_11 ? 2'h0 : _ctrl_T_409; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_411 = _ctrl_T_9 ? 2'h0 : _ctrl_T_410; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_412 = _ctrl_T_7 ? 2'h0 : _ctrl_T_411; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_413 = _ctrl_T_5 ? 2'h0 : _ctrl_T_412; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_414 = _ctrl_T_3 ? 2'h0 : _ctrl_T_413; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_433 = _ctrl_T_83 ? 2'h3 : _ctrl_T_373; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_434 = _ctrl_T_81 ? 2'h2 : _ctrl_T_433; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_435 = _ctrl_T_79 ? 2'h0 : _ctrl_T_434; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_436 = _ctrl_T_77 ? 2'h0 : _ctrl_T_435; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_437 = _ctrl_T_75 ? 2'h0 : _ctrl_T_436; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_438 = _ctrl_T_73 ? 2'h0 : _ctrl_T_437; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_439 = _ctrl_T_71 ? 2'h0 : _ctrl_T_438; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_440 = _ctrl_T_69 ? 2'h0 : _ctrl_T_439; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_441 = _ctrl_T_67 ? 2'h0 : _ctrl_T_440; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_442 = _ctrl_T_65 ? 2'h0 : _ctrl_T_441; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_443 = _ctrl_T_63 ? 2'h0 : _ctrl_T_442; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_444 = _ctrl_T_61 ? 2'h0 : _ctrl_T_443; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_445 = _ctrl_T_59 ? 2'h0 : _ctrl_T_444; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_446 = _ctrl_T_57 ? 2'h0 : _ctrl_T_445; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_447 = _ctrl_T_55 ? 2'h0 : _ctrl_T_446; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_448 = _ctrl_T_53 ? 2'h0 : _ctrl_T_447; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_449 = _ctrl_T_51 ? 2'h0 : _ctrl_T_448; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_450 = _ctrl_T_49 ? 2'h0 : _ctrl_T_449; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_451 = _ctrl_T_47 ? 2'h0 : _ctrl_T_450; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_452 = _ctrl_T_45 ? 2'h0 : _ctrl_T_451; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_453 = _ctrl_T_43 ? 2'h0 : _ctrl_T_452; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_454 = _ctrl_T_41 ? 2'h0 : _ctrl_T_453; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_455 = _ctrl_T_39 ? 2'h0 : _ctrl_T_454; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_456 = _ctrl_T_37 ? 2'h0 : _ctrl_T_455; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_457 = _ctrl_T_35 ? 2'h2 : _ctrl_T_456; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_458 = _ctrl_T_33 ? 2'h1 : _ctrl_T_457; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_459 = _ctrl_T_31 ? 2'h0 : _ctrl_T_458; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_460 = _ctrl_T_29 ? 2'h1 : _ctrl_T_459; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_461 = _ctrl_T_27 ? 2'h0 : _ctrl_T_460; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_462 = _ctrl_T_25 ? 2'h2 : _ctrl_T_461; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_463 = _ctrl_T_23 ? 2'h1 : _ctrl_T_462; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_464 = _ctrl_T_21 ? 2'h0 : _ctrl_T_463; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_465 = _ctrl_T_19 ? 2'h0 : _ctrl_T_464; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_466 = _ctrl_T_17 ? 2'h0 : _ctrl_T_465; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_467 = _ctrl_T_15 ? 2'h0 : _ctrl_T_466; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_468 = _ctrl_T_13 ? 2'h0 : _ctrl_T_467; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_469 = _ctrl_T_11 ? 2'h0 : _ctrl_T_468; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_470 = _ctrl_T_9 ? 2'h0 : _ctrl_T_469; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_471 = _ctrl_T_7 ? 2'h0 : _ctrl_T_470; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_472 = _ctrl_T_5 ? 2'h0 : _ctrl_T_471; // @[Lookup.scala 33:37]
  wire [1:0] _ctrl_T_473 = _ctrl_T_3 ? 2'h0 : _ctrl_T_472; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_476 = _ctrl_T_115 ? 3'h3 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_477 = _ctrl_T_113 ? 3'h2 : _ctrl_T_476; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_478 = _ctrl_T_111 ? 3'h1 : _ctrl_T_477; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_479 = _ctrl_T_109 ? 3'h3 : _ctrl_T_478; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_480 = _ctrl_T_107 ? 3'h2 : _ctrl_T_479; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_481 = _ctrl_T_105 ? 3'h1 : _ctrl_T_480; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_482 = _ctrl_T_103 ? 3'h0 : _ctrl_T_481; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_483 = _ctrl_T_101 ? 3'h0 : _ctrl_T_482; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_484 = _ctrl_T_99 ? 3'h0 : _ctrl_T_483; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_485 = _ctrl_T_97 ? 3'h0 : _ctrl_T_484; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_486 = _ctrl_T_95 ? 3'h0 : _ctrl_T_485; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_487 = _ctrl_T_93 ? 3'h0 : _ctrl_T_486; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_488 = _ctrl_T_91 ? 3'h0 : _ctrl_T_487; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_489 = _ctrl_T_89 ? 3'h0 : _ctrl_T_488; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_490 = _ctrl_T_87 ? 3'h0 : _ctrl_T_489; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_491 = _ctrl_T_85 ? 3'h0 : _ctrl_T_490; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_492 = _ctrl_T_83 ? 3'h0 : _ctrl_T_491; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_493 = _ctrl_T_81 ? 3'h0 : _ctrl_T_492; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_494 = _ctrl_T_79 ? 3'h0 : _ctrl_T_493; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_495 = _ctrl_T_77 ? 3'h5 : _ctrl_T_494; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_496 = _ctrl_T_75 ? 3'h4 : _ctrl_T_495; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_497 = _ctrl_T_73 ? 3'h0 : _ctrl_T_496; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_498 = _ctrl_T_71 ? 3'h0 : _ctrl_T_497; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_499 = _ctrl_T_69 ? 3'h0 : _ctrl_T_498; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_500 = _ctrl_T_67 ? 3'h0 : _ctrl_T_499; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_501 = _ctrl_T_65 ? 3'h0 : _ctrl_T_500; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_502 = _ctrl_T_63 ? 3'h0 : _ctrl_T_501; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_503 = _ctrl_T_61 ? 3'h0 : _ctrl_T_502; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_504 = _ctrl_T_59 ? 3'h0 : _ctrl_T_503; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_505 = _ctrl_T_57 ? 3'h0 : _ctrl_T_504; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_506 = _ctrl_T_55 ? 3'h0 : _ctrl_T_505; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_507 = _ctrl_T_53 ? 3'h0 : _ctrl_T_506; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_508 = _ctrl_T_51 ? 3'h0 : _ctrl_T_507; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_509 = _ctrl_T_49 ? 3'h0 : _ctrl_T_508; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_510 = _ctrl_T_47 ? 3'h0 : _ctrl_T_509; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_511 = _ctrl_T_45 ? 3'h0 : _ctrl_T_510; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_512 = _ctrl_T_43 ? 3'h0 : _ctrl_T_511; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_513 = _ctrl_T_41 ? 3'h0 : _ctrl_T_512; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_514 = _ctrl_T_39 ? 3'h0 : _ctrl_T_513; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_515 = _ctrl_T_37 ? 3'h0 : _ctrl_T_514; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_516 = _ctrl_T_35 ? 3'h0 : _ctrl_T_515; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_517 = _ctrl_T_33 ? 3'h0 : _ctrl_T_516; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_518 = _ctrl_T_31 ? 3'h0 : _ctrl_T_517; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_519 = _ctrl_T_29 ? 3'h0 : _ctrl_T_518; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_520 = _ctrl_T_27 ? 3'h0 : _ctrl_T_519; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_521 = _ctrl_T_25 ? 3'h0 : _ctrl_T_520; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_522 = _ctrl_T_23 ? 3'h0 : _ctrl_T_521; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_523 = _ctrl_T_21 ? 3'h0 : _ctrl_T_522; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_524 = _ctrl_T_19 ? 3'h0 : _ctrl_T_523; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_525 = _ctrl_T_17 ? 3'h0 : _ctrl_T_524; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_526 = _ctrl_T_15 ? 3'h0 : _ctrl_T_525; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_527 = _ctrl_T_13 ? 3'h0 : _ctrl_T_526; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_528 = _ctrl_T_11 ? 3'h0 : _ctrl_T_527; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_529 = _ctrl_T_9 ? 3'h0 : _ctrl_T_528; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_530 = _ctrl_T_7 ? 3'h0 : _ctrl_T_529; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_531 = _ctrl_T_5 ? 3'h0 : _ctrl_T_530; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_532 = _ctrl_T_3 ? 3'h0 : _ctrl_T_531; // @[Lookup.scala 33:37]
  wire  _ctrl_T_550 = _ctrl_T_85 ? 1'h0 : _ctrl_T_87 | (_ctrl_T_89 | (_ctrl_T_91 | (_ctrl_T_93 | (_ctrl_T_95 | (
    _ctrl_T_97 | (_ctrl_T_99 | (_ctrl_T_101 | _ctrl_T_103))))))); // @[Lookup.scala 33:37]
  wire  _ctrl_T_551 = _ctrl_T_83 ? 1'h0 : _ctrl_T_550; // @[Lookup.scala 33:37]
  wire  _ctrl_T_552 = _ctrl_T_81 ? 1'h0 : _ctrl_T_551; // @[Lookup.scala 33:37]
  wire  _ctrl_T_553 = _ctrl_T_79 ? 1'h0 : _ctrl_T_552; // @[Lookup.scala 33:37]
  wire  _ctrl_T_554 = _ctrl_T_77 ? 1'h0 : _ctrl_T_553; // @[Lookup.scala 33:37]
  wire  _ctrl_T_555 = _ctrl_T_75 ? 1'h0 : _ctrl_T_554; // @[Lookup.scala 33:37]
  wire  _ctrl_T_556 = _ctrl_T_73 ? 1'h0 : _ctrl_T_555; // @[Lookup.scala 33:37]
  wire  _ctrl_T_557 = _ctrl_T_71 ? 1'h0 : _ctrl_T_556; // @[Lookup.scala 33:37]
  wire  _ctrl_T_558 = _ctrl_T_69 ? 1'h0 : _ctrl_T_557; // @[Lookup.scala 33:37]
  wire  _ctrl_T_559 = _ctrl_T_67 ? 1'h0 : _ctrl_T_558; // @[Lookup.scala 33:37]
  wire  _ctrl_T_560 = _ctrl_T_65 ? 1'h0 : _ctrl_T_559; // @[Lookup.scala 33:37]
  wire  _ctrl_T_561 = _ctrl_T_63 ? 1'h0 : _ctrl_T_560; // @[Lookup.scala 33:37]
  wire  _ctrl_T_562 = _ctrl_T_61 ? 1'h0 : _ctrl_T_561; // @[Lookup.scala 33:37]
  wire  _ctrl_T_563 = _ctrl_T_59 ? 1'h0 : _ctrl_T_562; // @[Lookup.scala 33:37]
  wire  _ctrl_T_564 = _ctrl_T_57 ? 1'h0 : _ctrl_T_563; // @[Lookup.scala 33:37]
  wire  _ctrl_T_565 = _ctrl_T_55 ? 1'h0 : _ctrl_T_564; // @[Lookup.scala 33:37]
  wire  _ctrl_T_566 = _ctrl_T_53 ? 1'h0 : _ctrl_T_565; // @[Lookup.scala 33:37]
  wire  _ctrl_T_567 = _ctrl_T_51 ? 1'h0 : _ctrl_T_566; // @[Lookup.scala 33:37]
  wire  _ctrl_T_568 = _ctrl_T_49 ? 1'h0 : _ctrl_T_567; // @[Lookup.scala 33:37]
  wire  _ctrl_T_569 = _ctrl_T_47 ? 1'h0 : _ctrl_T_568; // @[Lookup.scala 33:37]
  wire  _ctrl_T_570 = _ctrl_T_45 ? 1'h0 : _ctrl_T_569; // @[Lookup.scala 33:37]
  wire  _ctrl_T_571 = _ctrl_T_43 ? 1'h0 : _ctrl_T_570; // @[Lookup.scala 33:37]
  wire  _ctrl_T_572 = _ctrl_T_41 ? 1'h0 : _ctrl_T_571; // @[Lookup.scala 33:37]
  wire  _ctrl_T_573 = _ctrl_T_39 ? 1'h0 : _ctrl_T_572; // @[Lookup.scala 33:37]
  wire  _ctrl_T_574 = _ctrl_T_37 ? 1'h0 : _ctrl_T_573; // @[Lookup.scala 33:37]
  wire  _ctrl_T_575 = _ctrl_T_35 ? 1'h0 : _ctrl_T_574; // @[Lookup.scala 33:37]
  wire  _ctrl_T_576 = _ctrl_T_33 ? 1'h0 : _ctrl_T_575; // @[Lookup.scala 33:37]
  wire  _ctrl_T_577 = _ctrl_T_31 ? 1'h0 : _ctrl_T_576; // @[Lookup.scala 33:37]
  wire  _ctrl_T_578 = _ctrl_T_29 ? 1'h0 : _ctrl_T_577; // @[Lookup.scala 33:37]
  wire  _ctrl_T_579 = _ctrl_T_27 ? 1'h0 : _ctrl_T_578; // @[Lookup.scala 33:37]
  wire  _ctrl_T_580 = _ctrl_T_25 ? 1'h0 : _ctrl_T_579; // @[Lookup.scala 33:37]
  wire  _ctrl_T_581 = _ctrl_T_23 ? 1'h0 : _ctrl_T_580; // @[Lookup.scala 33:37]
  wire  _ctrl_T_582 = _ctrl_T_21 ? 1'h0 : _ctrl_T_581; // @[Lookup.scala 33:37]
  wire  _ctrl_T_583 = _ctrl_T_19 ? 1'h0 : _ctrl_T_582; // @[Lookup.scala 33:37]
  wire  _ctrl_T_584 = _ctrl_T_17 ? 1'h0 : _ctrl_T_583; // @[Lookup.scala 33:37]
  wire  _ctrl_T_585 = _ctrl_T_15 ? 1'h0 : _ctrl_T_584; // @[Lookup.scala 33:37]
  wire  _ctrl_T_586 = _ctrl_T_13 ? 1'h0 : _ctrl_T_585; // @[Lookup.scala 33:37]
  wire  _ctrl_T_587 = _ctrl_T_11 ? 1'h0 : _ctrl_T_586; // @[Lookup.scala 33:37]
  wire  _ctrl_T_588 = _ctrl_T_9 ? 1'h0 : _ctrl_T_587; // @[Lookup.scala 33:37]
  wire  _ctrl_T_589 = _ctrl_T_7 ? 1'h0 : _ctrl_T_588; // @[Lookup.scala 33:37]
  wire  _ctrl_T_590 = _ctrl_T_5 ? 1'h0 : _ctrl_T_589; // @[Lookup.scala 33:37]
  wire  _ctrl_T_591 = _ctrl_T_3 ? 1'h0 : _ctrl_T_590; // @[Lookup.scala 33:37]
  wire  c0_0 = _ctrl_T_1 ? 1'h0 : _ctrl_T_591; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_594 = _ctrl_T_115 ? 3'h2 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_595 = _ctrl_T_113 ? 3'h2 : _ctrl_T_594; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_596 = _ctrl_T_111 ? 3'h2 : _ctrl_T_595; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_597 = _ctrl_T_109 ? 3'h1 : _ctrl_T_596; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_598 = _ctrl_T_107 ? 3'h1 : _ctrl_T_597; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_599 = _ctrl_T_105 ? 3'h1 : _ctrl_T_598; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_600 = _ctrl_T_103 ? 3'h1 : _ctrl_T_599; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_601 = _ctrl_T_101 ? 3'h1 : _ctrl_T_600; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_602 = _ctrl_T_99 ? 3'h1 : _ctrl_T_601; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_603 = _ctrl_T_97 ? 3'h1 : _ctrl_T_602; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_604 = _ctrl_T_95 ? 3'h1 : _ctrl_T_603; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_605 = _ctrl_T_93 ? 3'h1 : _ctrl_T_604; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_606 = _ctrl_T_91 ? 3'h1 : _ctrl_T_605; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_607 = _ctrl_T_89 ? 3'h1 : _ctrl_T_606; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_608 = _ctrl_T_87 ? 3'h1 : _ctrl_T_607; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_609 = _ctrl_T_85 ? 3'h1 : _ctrl_T_608; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_610 = _ctrl_T_83 ? 3'h1 : _ctrl_T_609; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_611 = _ctrl_T_81 ? 3'h1 : _ctrl_T_610; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_612 = _ctrl_T_79 ? 3'h0 : _ctrl_T_611; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_613 = _ctrl_T_77 ? 3'h0 : _ctrl_T_612; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_614 = _ctrl_T_75 ? 3'h0 : _ctrl_T_613; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_615 = _ctrl_T_73 ? 3'h1 : _ctrl_T_614; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_616 = _ctrl_T_71 ? 3'h1 : _ctrl_T_615; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_617 = _ctrl_T_69 ? 3'h1 : _ctrl_T_616; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_618 = _ctrl_T_67 ? 3'h1 : _ctrl_T_617; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_619 = _ctrl_T_65 ? 3'h1 : _ctrl_T_618; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_620 = _ctrl_T_63 ? 3'h1 : _ctrl_T_619; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_621 = _ctrl_T_61 ? 3'h1 : _ctrl_T_620; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_622 = _ctrl_T_59 ? 3'h1 : _ctrl_T_621; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_623 = _ctrl_T_57 ? 3'h1 : _ctrl_T_622; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_624 = _ctrl_T_55 ? 3'h1 : _ctrl_T_623; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_625 = _ctrl_T_53 ? 3'h1 : _ctrl_T_624; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_626 = _ctrl_T_51 ? 3'h1 : _ctrl_T_625; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_627 = _ctrl_T_49 ? 3'h1 : _ctrl_T_626; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_628 = _ctrl_T_47 ? 3'h1 : _ctrl_T_627; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_629 = _ctrl_T_45 ? 3'h1 : _ctrl_T_628; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_630 = _ctrl_T_43 ? 3'h1 : _ctrl_T_629; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_631 = _ctrl_T_41 ? 3'h1 : _ctrl_T_630; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_632 = _ctrl_T_39 ? 3'h1 : _ctrl_T_631; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_633 = _ctrl_T_37 ? 3'h1 : _ctrl_T_632; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_634 = _ctrl_T_35 ? 3'h1 : _ctrl_T_633; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_635 = _ctrl_T_33 ? 3'h1 : _ctrl_T_634; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_636 = _ctrl_T_31 ? 3'h1 : _ctrl_T_635; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_637 = _ctrl_T_29 ? 3'h1 : _ctrl_T_636; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_638 = _ctrl_T_27 ? 3'h1 : _ctrl_T_637; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_639 = _ctrl_T_25 ? 3'h1 : _ctrl_T_638; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_640 = _ctrl_T_23 ? 3'h1 : _ctrl_T_639; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_641 = _ctrl_T_21 ? 3'h1 : _ctrl_T_640; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_642 = _ctrl_T_19 ? 3'h1 : _ctrl_T_641; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_643 = _ctrl_T_17 ? 3'h1 : _ctrl_T_642; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_644 = _ctrl_T_15 ? 3'h1 : _ctrl_T_643; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_645 = _ctrl_T_13 ? 3'h1 : _ctrl_T_644; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_646 = _ctrl_T_11 ? 3'h1 : _ctrl_T_645; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_647 = _ctrl_T_9 ? 3'h1 : _ctrl_T_646; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_648 = _ctrl_T_7 ? 3'h1 : _ctrl_T_647; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_649 = _ctrl_T_5 ? 3'h4 : _ctrl_T_648; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_650 = _ctrl_T_3 ? 3'h4 : _ctrl_T_649; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_659 = _ctrl_T_103 ? 3'h1 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_660 = _ctrl_T_101 ? 3'h1 : _ctrl_T_659; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_661 = _ctrl_T_99 ? 3'h1 : _ctrl_T_660; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_662 = _ctrl_T_97 ? 3'h1 : _ctrl_T_661; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_663 = _ctrl_T_95 ? 3'h1 : _ctrl_T_662; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_664 = _ctrl_T_93 ? 3'h2 : _ctrl_T_663; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_665 = _ctrl_T_91 ? 3'h2 : _ctrl_T_664; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_666 = _ctrl_T_89 ? 3'h2 : _ctrl_T_665; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_667 = _ctrl_T_87 ? 3'h2 : _ctrl_T_666; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_668 = _ctrl_T_85 ? 3'h1 : _ctrl_T_667; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_669 = _ctrl_T_83 ? 3'h2 : _ctrl_T_668; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_670 = _ctrl_T_81 ? 3'h2 : _ctrl_T_669; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_671 = _ctrl_T_79 ? 3'h0 : _ctrl_T_670; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_672 = _ctrl_T_77 ? 3'h0 : _ctrl_T_671; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_673 = _ctrl_T_75 ? 3'h0 : _ctrl_T_672; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_674 = _ctrl_T_73 ? 3'h1 : _ctrl_T_673; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_675 = _ctrl_T_71 ? 3'h1 : _ctrl_T_674; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_676 = _ctrl_T_69 ? 3'h1 : _ctrl_T_675; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_677 = _ctrl_T_67 ? 3'h1 : _ctrl_T_676; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_678 = _ctrl_T_65 ? 3'h1 : _ctrl_T_677; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_679 = _ctrl_T_63 ? 3'h1 : _ctrl_T_678; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_680 = _ctrl_T_61 ? 3'h1 : _ctrl_T_679; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_681 = _ctrl_T_59 ? 3'h1 : _ctrl_T_680; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_682 = _ctrl_T_57 ? 3'h1 : _ctrl_T_681; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_683 = _ctrl_T_55 ? 3'h1 : _ctrl_T_682; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_684 = _ctrl_T_53 ? 3'h2 : _ctrl_T_683; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_685 = _ctrl_T_51 ? 3'h2 : _ctrl_T_684; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_686 = _ctrl_T_49 ? 3'h2 : _ctrl_T_685; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_687 = _ctrl_T_47 ? 3'h2 : _ctrl_T_686; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_688 = _ctrl_T_45 ? 3'h2 : _ctrl_T_687; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_689 = _ctrl_T_43 ? 3'h2 : _ctrl_T_688; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_690 = _ctrl_T_41 ? 3'h2 : _ctrl_T_689; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_691 = _ctrl_T_39 ? 3'h2 : _ctrl_T_690; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_692 = _ctrl_T_37 ? 3'h2 : _ctrl_T_691; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_693 = _ctrl_T_35 ? 3'h1 : _ctrl_T_692; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_694 = _ctrl_T_33 ? 3'h1 : _ctrl_T_693; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_695 = _ctrl_T_31 ? 3'h1 : _ctrl_T_694; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_696 = _ctrl_T_29 ? 3'h2 : _ctrl_T_695; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_697 = _ctrl_T_27 ? 3'h2 : _ctrl_T_696; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_698 = _ctrl_T_25 ? 3'h2 : _ctrl_T_697; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_699 = _ctrl_T_23 ? 3'h2 : _ctrl_T_698; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_700 = _ctrl_T_21 ? 3'h2 : _ctrl_T_699; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_701 = _ctrl_T_19 ? 3'h1 : _ctrl_T_700; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_702 = _ctrl_T_17 ? 3'h1 : _ctrl_T_701; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_703 = _ctrl_T_15 ? 3'h1 : _ctrl_T_702; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_704 = _ctrl_T_13 ? 3'h1 : _ctrl_T_703; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_705 = _ctrl_T_11 ? 3'h1 : _ctrl_T_704; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_706 = _ctrl_T_9 ? 3'h1 : _ctrl_T_705; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_707 = _ctrl_T_7 ? 3'h1 : _ctrl_T_706; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_708 = _ctrl_T_5 ? 3'h2 : _ctrl_T_707; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_709 = _ctrl_T_3 ? 3'h2 : _ctrl_T_708; // @[Lookup.scala 33:37]
  wire  _ctrl_T_727 = _ctrl_T_85 ? 1'h0 : _ctrl_T_87 | (_ctrl_T_89 | (_ctrl_T_91 | (_ctrl_T_93 | (_ctrl_T_95 | (
    _ctrl_T_97 | (_ctrl_T_99 | (_ctrl_T_101 | (_ctrl_T_103 | (_ctrl_T_105 | (_ctrl_T_107 | (_ctrl_T_109 | (_ctrl_T_111
     | (_ctrl_T_113 | _ctrl_T_115))))))))))))); // @[Lookup.scala 33:37]
  wire  _ctrl_T_730 = _ctrl_T_79 ? 1'h0 : _ctrl_T_81 | (_ctrl_T_83 | _ctrl_T_727); // @[Lookup.scala 33:37]
  wire  _ctrl_T_731 = _ctrl_T_77 ? 1'h0 : _ctrl_T_730; // @[Lookup.scala 33:37]
  wire  _ctrl_T_732 = _ctrl_T_75 ? 1'h0 : _ctrl_T_731; // @[Lookup.scala 33:37]
  wire  _ctrl_T_752 = _ctrl_T_35 ? 1'h0 : _ctrl_T_37 | (_ctrl_T_39 | (_ctrl_T_41 | (_ctrl_T_43 | (_ctrl_T_45 | (
    _ctrl_T_47 | (_ctrl_T_49 | (_ctrl_T_51 | (_ctrl_T_53 | (_ctrl_T_55 | (_ctrl_T_57 | (_ctrl_T_59 | (_ctrl_T_61 | (
    _ctrl_T_63 | (_ctrl_T_65 | (_ctrl_T_67 | (_ctrl_T_69 | (_ctrl_T_71 | (_ctrl_T_73 | _ctrl_T_732)))))))))))))))))); // @[Lookup.scala 33:37]
  wire  _ctrl_T_753 = _ctrl_T_33 ? 1'h0 : _ctrl_T_752; // @[Lookup.scala 33:37]
  wire  _ctrl_T_754 = _ctrl_T_31 ? 1'h0 : _ctrl_T_753; // @[Lookup.scala 33:37]
  wire  _ctrl_T_760 = _ctrl_T_19 ? 1'h0 : _ctrl_T_21 | (_ctrl_T_23 | (_ctrl_T_25 | (_ctrl_T_27 | (_ctrl_T_29 |
    _ctrl_T_754)))); // @[Lookup.scala 33:37]
  wire  _ctrl_T_761 = _ctrl_T_17 ? 1'h0 : _ctrl_T_760; // @[Lookup.scala 33:37]
  wire  _ctrl_T_762 = _ctrl_T_15 ? 1'h0 : _ctrl_T_761; // @[Lookup.scala 33:37]
  wire  _ctrl_T_763 = _ctrl_T_13 ? 1'h0 : _ctrl_T_762; // @[Lookup.scala 33:37]
  wire  _ctrl_T_764 = _ctrl_T_11 ? 1'h0 : _ctrl_T_763; // @[Lookup.scala 33:37]
  wire  _ctrl_T_765 = _ctrl_T_9 ? 1'h0 : _ctrl_T_764; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_771 = _ctrl_T_115 ? 3'h7 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_772 = _ctrl_T_113 ? 3'h7 : _ctrl_T_771; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_773 = _ctrl_T_111 ? 3'h7 : _ctrl_T_772; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_774 = _ctrl_T_109 ? 3'h0 : _ctrl_T_773; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_775 = _ctrl_T_107 ? 3'h0 : _ctrl_T_774; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_776 = _ctrl_T_105 ? 3'h0 : _ctrl_T_775; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_777 = _ctrl_T_103 ? 3'h0 : _ctrl_T_776; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_778 = _ctrl_T_101 ? 3'h0 : _ctrl_T_777; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_779 = _ctrl_T_99 ? 3'h0 : _ctrl_T_778; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_780 = _ctrl_T_97 ? 3'h0 : _ctrl_T_779; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_781 = _ctrl_T_95 ? 3'h0 : _ctrl_T_780; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_782 = _ctrl_T_93 ? 3'h1 : _ctrl_T_781; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_783 = _ctrl_T_91 ? 3'h1 : _ctrl_T_782; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_784 = _ctrl_T_89 ? 3'h1 : _ctrl_T_783; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_785 = _ctrl_T_87 ? 3'h1 : _ctrl_T_784; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_786 = _ctrl_T_85 ? 3'h2 : _ctrl_T_785; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_787 = _ctrl_T_83 ? 3'h1 : _ctrl_T_786; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_788 = _ctrl_T_81 ? 3'h1 : _ctrl_T_787; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_789 = _ctrl_T_79 ? 3'h0 : _ctrl_T_788; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_790 = _ctrl_T_77 ? 3'h0 : _ctrl_T_789; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_791 = _ctrl_T_75 ? 3'h0 : _ctrl_T_790; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_792 = _ctrl_T_73 ? 3'h0 : _ctrl_T_791; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_793 = _ctrl_T_71 ? 3'h0 : _ctrl_T_792; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_794 = _ctrl_T_69 ? 3'h0 : _ctrl_T_793; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_795 = _ctrl_T_67 ? 3'h0 : _ctrl_T_794; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_796 = _ctrl_T_65 ? 3'h0 : _ctrl_T_795; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_797 = _ctrl_T_63 ? 3'h0 : _ctrl_T_796; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_798 = _ctrl_T_61 ? 3'h0 : _ctrl_T_797; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_799 = _ctrl_T_59 ? 3'h0 : _ctrl_T_798; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_800 = _ctrl_T_57 ? 3'h0 : _ctrl_T_799; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_801 = _ctrl_T_55 ? 3'h0 : _ctrl_T_800; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_802 = _ctrl_T_53 ? 3'h6 : _ctrl_T_801; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_803 = _ctrl_T_51 ? 3'h6 : _ctrl_T_802; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_804 = _ctrl_T_49 ? 3'h6 : _ctrl_T_803; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_805 = _ctrl_T_47 ? 3'h1 : _ctrl_T_804; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_806 = _ctrl_T_45 ? 3'h1 : _ctrl_T_805; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_807 = _ctrl_T_43 ? 3'h1 : _ctrl_T_806; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_808 = _ctrl_T_41 ? 3'h1 : _ctrl_T_807; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_809 = _ctrl_T_39 ? 3'h1 : _ctrl_T_808; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_810 = _ctrl_T_37 ? 3'h1 : _ctrl_T_809; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_811 = _ctrl_T_35 ? 3'h2 : _ctrl_T_810; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_812 = _ctrl_T_33 ? 3'h2 : _ctrl_T_811; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_813 = _ctrl_T_31 ? 3'h2 : _ctrl_T_812; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_814 = _ctrl_T_29 ? 3'h1 : _ctrl_T_813; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_815 = _ctrl_T_27 ? 3'h1 : _ctrl_T_814; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_816 = _ctrl_T_25 ? 3'h1 : _ctrl_T_815; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_817 = _ctrl_T_23 ? 3'h1 : _ctrl_T_816; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_818 = _ctrl_T_21 ? 3'h1 : _ctrl_T_817; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_819 = _ctrl_T_19 ? 3'h3 : _ctrl_T_818; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_820 = _ctrl_T_17 ? 3'h3 : _ctrl_T_819; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_821 = _ctrl_T_15 ? 3'h3 : _ctrl_T_820; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_822 = _ctrl_T_13 ? 3'h3 : _ctrl_T_821; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_823 = _ctrl_T_11 ? 3'h3 : _ctrl_T_822; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_824 = _ctrl_T_9 ? 3'h3 : _ctrl_T_823; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_825 = _ctrl_T_7 ? 3'h1 : _ctrl_T_824; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_826 = _ctrl_T_5 ? 3'h5 : _ctrl_T_825; // @[Lookup.scala 33:37]
  wire [2:0] _ctrl_T_827 = _ctrl_T_3 ? 3'h4 : _ctrl_T_826; // @[Lookup.scala 33:37]
  wire [2:0] c0_4 = _ctrl_T_1 ? 3'h4 : _ctrl_T_827; // @[Lookup.scala 33:37]
  wire [20:0] imm_i_hi = inst[31] ? 21'h1fffff : 21'h0; // @[Bitwise.scala 72:12]
  wire [10:0] imm_i_lo = inst[30:20]; // @[Decode.scala 117:43]
  wire [31:0] imm_i = {imm_i_hi,imm_i_lo}; // @[Cat.scala 30:58]
  wire [5:0] imm_s_hi_lo = inst[30:25]; // @[Decode.scala 118:43]
  wire [31:0] imm_s = {imm_i_hi,imm_s_hi_lo,inst[11:7]}; // @[Cat.scala 30:58]
  wire [19:0] imm_b_hi_hi_hi = inst[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire  imm_b_hi_hi_lo = inst[7]; // @[Decode.scala 119:43]
  wire [3:0] imm_b_lo_hi = inst[11:8]; // @[Decode.scala 119:66]
  wire [31:0] imm_b = {imm_b_hi_hi_hi,imm_b_hi_hi_lo,imm_s_hi_lo,imm_b_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [19:0] imm_u_hi = inst[31:12]; // @[Decode.scala 120:23]
  wire [31:0] imm_u = {imm_u_hi,12'h0}; // @[Cat.scala 30:58]
  wire [11:0] imm_j_hi_hi_hi = inst[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [7:0] imm_j_hi_hi_lo = inst[19:12]; // @[Decode.scala 121:43]
  wire  imm_j_hi_lo = inst[20]; // @[Decode.scala 121:57]
  wire [9:0] imm_j_lo_hi = inst[30:21]; // @[Decode.scala 121:67]
  wire [31:0] imm_j = {imm_j_hi_hi_hi,imm_j_hi_hi_lo,imm_j_hi_lo,imm_j_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [31:0] _imm_shamt_T = {27'h0,inst[24:20]}; // @[Cat.scala 30:58]
  wire [5:0] imm_shamt_lo_1 = inst[25:20]; // @[Decode.scala 122:88]
  wire [31:0] _imm_shamt_T_1 = {26'h0,imm_shamt_lo_1}; // @[Cat.scala 30:58]
  wire [31:0] imm_shamt = c0_0 ? _imm_shamt_T : _imm_shamt_T_1; // @[Decode.scala 122:22]
  wire [31:0] imm_csr = {27'h0,inst[19:15]}; // @[Cat.scala 30:58]
  wire [31:0] _io_out_bits_imm_T_1 = 3'h1 == c0_4 ? imm_i : 32'h0; // @[Mux.scala 80:57]
  wire [31:0] _io_out_bits_imm_T_3 = 3'h2 == c0_4 ? imm_s : _io_out_bits_imm_T_1; // @[Mux.scala 80:57]
  wire [31:0] _io_out_bits_imm_T_5 = 3'h3 == c0_4 ? imm_b : _io_out_bits_imm_T_3; // @[Mux.scala 80:57]
  wire [31:0] _io_out_bits_imm_T_7 = 3'h4 == c0_4 ? imm_u : _io_out_bits_imm_T_5; // @[Mux.scala 80:57]
  wire [31:0] _io_out_bits_imm_T_9 = 3'h5 == c0_4 ? imm_j : _io_out_bits_imm_T_7; // @[Mux.scala 80:57]
  wire [31:0] _io_out_bits_imm_T_11 = 3'h6 == c0_4 ? imm_shamt : _io_out_bits_imm_T_9; // @[Mux.scala 80:57]
  wire  _stall_T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  stall = ~_stall_T; // @[Decode.scala 135:15]
  assign io_in_ready = ~stall; // @[Decode.scala 136:18]
  assign io_out_valid = 1'h1; // @[Decode.scala 137:16]
  assign io_out_bits_valid = io_in_bits_inst_valid; // @[Decode.scala 102:26]
  assign io_out_bits_pc = io_in_bits_pc; // @[Decode.scala 100:23]
  assign io_out_bits_inst = io_in_bits_inst; // @[Decode.scala 101:23]
  assign io_out_bits_fu_code = _ctrl_T_1 ? 3'h1 : _ctrl_T_237; // @[Lookup.scala 33:37]
  assign io_out_bits_alu_code = _ctrl_T_1 ? 4'h1 : _ctrl_T_296; // @[Lookup.scala 33:37]
  assign io_out_bits_jmp_code = _ctrl_T_1 ? 4'h0 : _ctrl_T_355; // @[Lookup.scala 33:37]
  assign io_out_bits_mem_code = _ctrl_T_1 ? 2'h0 : _ctrl_T_414; // @[Lookup.scala 33:37]
  assign io_out_bits_mem_size = _ctrl_T_1 ? 2'h0 : _ctrl_T_473; // @[Lookup.scala 33:37]
  assign io_out_bits_csr_code = _ctrl_T_1 ? 3'h0 : _ctrl_T_532; // @[Lookup.scala 33:37]
  assign io_out_bits_w_type = _ctrl_T_1 ? 1'h0 : _ctrl_T_591; // @[Lookup.scala 33:37]
  assign io_out_bits_rs1_src = _ctrl_T_1 ? 3'h3 : _ctrl_T_650; // @[Lookup.scala 33:37]
  assign io_out_bits_rs2_src = _ctrl_T_1 ? 3'h2 : _ctrl_T_709; // @[Lookup.scala 33:37]
  assign io_out_bits_rs1_addr = inst[19:15]; // @[Decode.scala 113:31]
  assign io_out_bits_rs2_addr = inst[24:20]; // @[Decode.scala 114:31]
  assign io_out_bits_rd_addr = inst[11:7]; // @[Decode.scala 115:30]
  assign io_out_bits_rd_en = _ctrl_T_1 | (_ctrl_T_3 | (_ctrl_T_5 | (_ctrl_T_7 | _ctrl_T_765))); // @[Lookup.scala 33:37]
  assign io_out_bits_imm = 3'h7 == c0_4 ? imm_csr : _io_out_bits_imm_T_11; // @[Mux.scala 80:57]
  always @(posedge clock) begin
    if (reset) begin // @[Decode.scala 15:22]
      inst <= 32'h0; // @[Decode.scala 15:22]
    end else if (_T) begin // @[Decode.scala 18:21]
      if (io_id_flush) begin // @[Decode.scala 20:16]
        inst <= 32'h0;
      end else begin
        inst <= io_in_bits_inst;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
